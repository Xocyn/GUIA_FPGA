architecture behavior of ejcombtb is 
component ejcomb
port (
		A: in std_logic;
		B: in std_logic;
		LED: out std_logic);
end component;

--inputs
signal A:std_logic:='0';
signal B:std_logic:='0';
--ouputs
signal LED:std_logic;

begin
--instantiate the units under test (uut)
uut: ejcomb port map (A=> A, B=> B, LED=> LED);

stimproc: process
begin
A<='0';B<='0'; wait for 10ns;
A<='0';B<='1'; wait for 10ns;
A<='1';B<='0'; wait for 10ns;
A<='1';B<='1'; wait for 10ns;
wait; 
end process;
end;
